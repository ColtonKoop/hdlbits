module top_module ( input a, input b, output out );
	
    mod_a mod_a1( a, b, out);
    
endmodule